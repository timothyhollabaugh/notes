library verilog;
use verilog.vl_types.all;
entity single_cycle_CPU_tb is
end single_cycle_CPU_tb;
