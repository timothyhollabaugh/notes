library verilog;
use verilog.vl_types.all;
entity lab_1_testbench is
end lab_1_testbench;
