
module Toplevel(CLOCK_50, SW, VGA_R, VGA_G, VGA_HS, VGA_VS, LEDG);
    input CLOCK_50;
    input [9:0] SW;
    output [9:0] LEDG;
    output [3:0] VGA_R, VGA_G;
    output VGA_HS, VGA_VS;

    wire [1200:0] data;

    wire [39:0] ctrl;

    assign ctrl = {SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0], SW[0]};


    assign data[  39:   0] = 40'b1111111111111111111111111111111111111111 ^ ctrl;
    assign data[  79:  40] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 119:  80] = 40'b1000000000000000000111000100010111010101 ^ ctrl;
    assign data[ 159: 120] = 40'b1000000000000000000101000100010001010101 ^ ctrl;
    assign data[ 199: 160] = 40'b1000000000000000000101000100010111011101 ^ ctrl;
    assign data[ 239: 200] = 40'b1000000000000000000101000100010001010101 ^ ctrl;
    assign data[ 279: 240] = 40'b1000000000000000010111011101110111010101 ^ ctrl;
    assign data[ 319: 280] = 40'b1000000000000000001000000000000000000001 ^ ctrl;
    assign data[ 359: 320] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 399: 360] = 40'b1000000000000001001100010011011101000101 ^ ctrl;
    assign data[ 439: 400] = 40'b1000000000000001010100010101010101000101 ^ ctrl;
    assign data[ 479: 440] = 40'b1000000000000001010100010011010101000101 ^ ctrl;
    assign data[ 519: 480] = 40'b1000000000000000010100010101010101010101 ^ ctrl;
    assign data[ 559: 520] = 40'b1000000000000001001101110101011100101001 ^ ctrl;
    assign data[ 599: 560] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 639: 600] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 679: 640] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 719: 680] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 759: 720] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 799: 760] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 839: 800] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 879: 840] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 919: 880] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 959: 920] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[ 999: 960] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[1039:1000] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[1079:1040] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[1119:1080] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[1159:1120] = 40'b1000000000000000000000000000000000000001 ^ ctrl;
    assign data[1199:1160] = 40'b1111111111111111111111111111111111111111 ^ ctrl;

    wire pixel_position;

    VGA_Test vga (
        .clk(CLOCK_50),
        .data(data),
        .red_out(VGA_R),
        .green_out(VGA_G),
        .h_sync_out(VGA_HS),
        .v_sync_out(VGA_VS),
    );

endmodule

